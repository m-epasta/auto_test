module main

fn test_add() {
    // TODO: Implement test for add
    assert true
}

